module Assets/snakeBody_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=10'b0000000000) && ({row_reg, col_reg}<10'b0000001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b0000001000) && ({row_reg, col_reg}<10'b0000001010)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0000001010)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0000001011)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0000001100) && ({row_reg, col_reg}<10'b0000001110)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0000001110)) color_data = 12'b100010010001;
		if(({row_reg, col_reg}>=10'b0000001111) && ({row_reg, col_reg}<10'b0000010001)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b0000010001)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0000010010)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0000010011)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0000010100)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0000010101)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b0000010110)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}>=10'b0000010111) && ({row_reg, col_reg}<10'b0000011001)) color_data = 12'b101111010001;

		if(({row_reg, col_reg}>=10'b0000011001) && ({row_reg, col_reg}<10'b0000100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==10'b0000100101)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0000100110) && ({row_reg, col_reg}<10'b0000101011)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0000101011)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0000101100) && ({row_reg, col_reg}<10'b0000101110)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0000101110)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b0000101111) && ({row_reg, col_reg}<10'b0000110001)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b0000110001)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0000110010) && ({row_reg, col_reg}<10'b0000110101)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0000110101)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0000110110)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0000110111)) color_data = 12'b101111110000;
		if(({row_reg, col_reg}>=10'b0000111000) && ({row_reg, col_reg}<10'b0000111011)) color_data = 12'b101111010001;

		if(({row_reg, col_reg}>=10'b0000111011) && ({row_reg, col_reg}<10'b0001000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b0001000010) && ({row_reg, col_reg}<10'b0001000101)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b0001000101) && ({row_reg, col_reg}<10'b0001000111)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0001000111)) color_data = 12'b101111100001;
		if(({row_reg, col_reg}>=10'b0001001000) && ({row_reg, col_reg}<10'b0001001010)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0001001010)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0001001011)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0001001100)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0001001101) && ({row_reg, col_reg}<10'b0001001111)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0001001111)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}>=10'b0001010000) && ({row_reg, col_reg}<10'b0001010010)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0001010010)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0001010011)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0001010100) && ({row_reg, col_reg}<10'b0001010110)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}>=10'b0001010110) && ({row_reg, col_reg}<10'b0001011000)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0001011000)) color_data = 12'b110011100001;
		if(({row_reg, col_reg}==10'b0001011001)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0001011010)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0001011011) && ({row_reg, col_reg}<10'b0001011101)) color_data = 12'b101010110001;

		if(({row_reg, col_reg}==10'b0001011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b0001100000) && ({row_reg, col_reg}<10'b0001100100)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0001100100)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b0001100101) && ({row_reg, col_reg}<10'b0001101000)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0001101000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0001101001)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0001101010)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}>=10'b0001101011) && ({row_reg, col_reg}<10'b0001101110)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0001101110)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0001101111)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0001110000) && ({row_reg, col_reg}<10'b0001110010)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}>=10'b0001110010) && ({row_reg, col_reg}<10'b0001110100)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}>=10'b0001110100) && ({row_reg, col_reg}<10'b0001111001)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0001111001)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0001111010)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0001111011)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0001111100)) color_data = 12'b011110010000;

		if(({row_reg, col_reg}==10'b0001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b0010000000) && ({row_reg, col_reg}<10'b0010000010)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b0010000010)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0010000011)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0010000100)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b0010000101)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b0010000110) && ({row_reg, col_reg}<10'b0010001000)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0010001000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0010001001)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}>=10'b0010001010) && ({row_reg, col_reg}<10'b0010001101)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0010001101) && ({row_reg, col_reg}<10'b0010001111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}>=10'b0010001111) && ({row_reg, col_reg}<10'b0010010011)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}>=10'b0010010011) && ({row_reg, col_reg}<10'b0010010101)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0010010101)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}>=10'b0010010110) && ({row_reg, col_reg}<10'b0010011000)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0010011000) && ({row_reg, col_reg}<10'b0010011010)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0010011010)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b0010011011) && ({row_reg, col_reg}<10'b0010011101)) color_data = 12'b100010100000;

		if(({row_reg, col_reg}==10'b0010011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b0010100000) && ({row_reg, col_reg}<10'b0010100010)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0010100010)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0010100011)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0010100100)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b0010100101) && ({row_reg, col_reg}<10'b0010101010)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0010101010)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0010101011)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}>=10'b0010101100) && ({row_reg, col_reg}<10'b0010101110)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}>=10'b0010101110) && ({row_reg, col_reg}<10'b0010110000)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}>=10'b0010110000) && ({row_reg, col_reg}<10'b0010110100)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0010110100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0010110101)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}>=10'b0010110110) && ({row_reg, col_reg}<10'b0010111000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0010111000)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0010111001)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0010111010) && ({row_reg, col_reg}<10'b0010111101)) color_data = 12'b100010100000;

		if(({row_reg, col_reg}==10'b0010111101)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0011000000) && ({row_reg, col_reg}<10'b0011000011)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0011000011)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0011000100)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0011000101)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0011000110) && ({row_reg, col_reg}<10'b0011001000)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0011001000)) color_data = 12'b110011100001;
		if(({row_reg, col_reg}==10'b0011001001)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}==10'b0011001010)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}>=10'b0011001011) && ({row_reg, col_reg}<10'b0011001101)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}>=10'b0011001101) && ({row_reg, col_reg}<10'b0011001111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0011001111)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0011010000)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0011010001) && ({row_reg, col_reg}<10'b0011010011)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0011010011)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0011010100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0011010101)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0011010110)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b0011010111)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0011011000)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}>=10'b0011011001) && ({row_reg, col_reg}<10'b0011011100)) color_data = 12'b100010010000;

		if(({row_reg, col_reg}>=10'b0011011100) && ({row_reg, col_reg}<10'b0011100011)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0011100011)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0011100100)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}>=10'b0011100101) && ({row_reg, col_reg}<10'b0011100111)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0011100111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0011101000)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}>=10'b0011101001) && ({row_reg, col_reg}<10'b0011101011)) color_data = 12'b110011100001;
		if(({row_reg, col_reg}==10'b0011101011)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0011101100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0011101101) && ({row_reg, col_reg}<10'b0011101111)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}>=10'b0011101111) && ({row_reg, col_reg}<10'b0011110001)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0011110001)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b0011110010) && ({row_reg, col_reg}<10'b0011110100)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b0011110100)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0011110101) && ({row_reg, col_reg}<10'b0011110111)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0011110111)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0011111000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0011111001)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0011111010)) color_data = 12'b100010010000;

		if(({row_reg, col_reg}>=10'b0011111011) && ({row_reg, col_reg}<10'b0100000000)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}>=10'b0100000000) && ({row_reg, col_reg}<10'b0100000100)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0100000100)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}>=10'b0100000101) && ({row_reg, col_reg}<10'b0100000111)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}>=10'b0100000111) && ({row_reg, col_reg}<10'b0100001001)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0100001001)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0100001010)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0100001011)) color_data = 12'b101011000000;
		if(({row_reg, col_reg}==10'b0100001100)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0100001101)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b0100001110) && ({row_reg, col_reg}<10'b0100010001)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0100010001) && ({row_reg, col_reg}<10'b0100010011)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}>=10'b0100010011) && ({row_reg, col_reg}<10'b0100010110)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0100010110) && ({row_reg, col_reg}<10'b0100011000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b0100011000) && ({row_reg, col_reg}<10'b0100011010)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b0100011010) && ({row_reg, col_reg}<10'b0100011101)) color_data = 12'b100010100000;

		if(({row_reg, col_reg}==10'b0100011101)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0100100000) && ({row_reg, col_reg}<10'b0100100010)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0100100010)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0100100011)) color_data = 12'b101011000000;
		if(({row_reg, col_reg}==10'b0100100100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0100100101)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0100100110)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0100100111)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0100101000)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0100101001)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}>=10'b0100101010) && ({row_reg, col_reg}<10'b0100101100)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0100101100)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0100101101)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b0100101110) && ({row_reg, col_reg}<10'b0100110000)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0100110000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b0100110001) && ({row_reg, col_reg}<10'b0100110100)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0100110100)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0100110101)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b0100110110) && ({row_reg, col_reg}<10'b0100111010)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0100111010) && ({row_reg, col_reg}<10'b0100111100)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0100111100)) color_data = 12'b100010010000;

		if(({row_reg, col_reg}==10'b0100111101)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0101000000)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0101000001) && ({row_reg, col_reg}<10'b0101000011)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0101000011)) color_data = 12'b101011000000;
		if(({row_reg, col_reg}==10'b0101000100)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0101000101)) color_data = 12'b110011100001;
		if(({row_reg, col_reg}==10'b0101000110)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0101000111)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}>=10'b0101001000) && ({row_reg, col_reg}<10'b0101001010)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0101001010)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0101001011) && ({row_reg, col_reg}<10'b0101001101)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0101001101)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0101001110) && ({row_reg, col_reg}<10'b0101010110)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b0101010110) && ({row_reg, col_reg}<10'b0101011001)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0101011001) && ({row_reg, col_reg}<10'b0101011101)) color_data = 12'b011110010000;

		if(({row_reg, col_reg}==10'b0101011101)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b0101100000) && ({row_reg, col_reg}<10'b0101100011)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0101100011)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0101100100)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}>=10'b0101100101) && ({row_reg, col_reg}<10'b0101100111)) color_data = 12'b110011100001;
		if(({row_reg, col_reg}==10'b0101100111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0101101000)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}>=10'b0101101001) && ({row_reg, col_reg}<10'b0101101011)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0101101011)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b0101101100) && ({row_reg, col_reg}<10'b0101101110)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b0101101110) && ({row_reg, col_reg}<10'b0101110010)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b0101110010) && ({row_reg, col_reg}<10'b0101110101)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0101110101)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0101110110)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0101110111)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0101111000)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0101111001)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b0101111010) && ({row_reg, col_reg}<10'b0101111101)) color_data = 12'b011110000000;

		if(({row_reg, col_reg}==10'b0101111101)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}>=10'b0110000000) && ({row_reg, col_reg}<10'b0110000011)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b0110000011)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0110000100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b0110000101) && ({row_reg, col_reg}<10'b0110000111)) color_data = 12'b110011100001;
		if(({row_reg, col_reg}==10'b0110000111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0110001000)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0110001001)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0110001010)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b0110001011) && ({row_reg, col_reg}<10'b0110010011)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0110010011)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0110010100)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0110010101) && ({row_reg, col_reg}<10'b0110011000)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0110011000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0110011001)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b0110011010) && ({row_reg, col_reg}<10'b0110011101)) color_data = 12'b010101100000;

		if(({row_reg, col_reg}==10'b0110011101)) color_data = 12'b010101010000;
		if(({row_reg, col_reg}>=10'b0110100000) && ({row_reg, col_reg}<10'b0110100011)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b0110100011)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b0110100100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0110100101)) color_data = 12'b110011100001;
		if(({row_reg, col_reg}>=10'b0110100110) && ({row_reg, col_reg}<10'b0110101000)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0110101000)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0110101001)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0110101010)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b0110101011) && ({row_reg, col_reg}<10'b0110101101)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0110101101)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b0110101110) && ({row_reg, col_reg}<10'b0110110011)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0110110011)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b0110110100) && ({row_reg, col_reg}<10'b0110110110)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b0110110110) && ({row_reg, col_reg}<10'b0110111000)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0110111000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b0110111001)) color_data = 12'b010101010000;

		if(({row_reg, col_reg}>=10'b0110111010) && ({row_reg, col_reg}<10'b0111000000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}>=10'b0111000000) && ({row_reg, col_reg}<10'b0111000011)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b0111000011)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0111000100)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0111000101)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}==10'b0111000110)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0111000111)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0111001000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0111001001)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}>=10'b0111001010) && ({row_reg, col_reg}<10'b0111001100)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0111001100)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0111001101)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0111001110)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0111001111)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0111010000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0111010001)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b0111010010)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b0111010011)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b0111010100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b0111010101)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b0111010110)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0111010111)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0111011000)) color_data = 12'b011001110000;

		if(({row_reg, col_reg}>=10'b0111011001) && ({row_reg, col_reg}<10'b0111100000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}>=10'b0111100000) && ({row_reg, col_reg}<10'b0111100011)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b0111100011)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b0111100100)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}>=10'b0111100101) && ({row_reg, col_reg}<10'b0111100111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b0111100111)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b0111101000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b0111101001)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b0111101010)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0111101011)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0111101100)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b0111101101)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b0111101110)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b0111101111)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0111110000)) color_data = 12'b011001100000;
		if(({row_reg, col_reg}==10'b0111110001)) color_data = 12'b001101000000;
		if(({row_reg, col_reg}>=10'b0111110010) && ({row_reg, col_reg}<10'b0111110100)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}==10'b0111110100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b0111110101) && ({row_reg, col_reg}<10'b0111110111)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b0111110111)) color_data = 12'b011001110000;

		if(({row_reg, col_reg}>=10'b0111111000) && ({row_reg, col_reg}<10'b1000000000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}>=10'b1000000000) && ({row_reg, col_reg}<10'b1000000011)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b1000000011)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b1000000100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1000000101)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1000000110)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}==10'b1000000111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1000001000)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b1000001001)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b1000001010)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}>=10'b1000001011) && ({row_reg, col_reg}<10'b1000001101)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b1000001101) && ({row_reg, col_reg}<10'b1000001111)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b1000001111)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1000010000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1000010001)) color_data = 12'b001101000000;
		if(({row_reg, col_reg}>=10'b1000010010) && ({row_reg, col_reg}<10'b1000010100)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}==10'b1000010100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1000010101)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b1000010110)) color_data = 12'b011001110000;

		if(({row_reg, col_reg}>=10'b1000010111) && ({row_reg, col_reg}<10'b1000100000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1000100000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b1000100001)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b1000100010)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b1000100011)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b1000100100)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b1000100101)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}>=10'b1000100110) && ({row_reg, col_reg}<10'b1000101000)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1000101000)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1000101001)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b1000101010)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b1000101011) && ({row_reg, col_reg}<10'b1000101101)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1000101101)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b1000101110) && ({row_reg, col_reg}<10'b1000110000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1000110000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1000110001)) color_data = 12'b001101000000;
		if(({row_reg, col_reg}>=10'b1000110010) && ({row_reg, col_reg}<10'b1000110100)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}==10'b1000110100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1000110101)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b1000110110)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1000110111)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1000111000)) color_data = 12'b010101110000;

		if(({row_reg, col_reg}>=10'b1000111001) && ({row_reg, col_reg}<10'b1001000000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}>=10'b1001000000) && ({row_reg, col_reg}<10'b1001000011)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b1001000011)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}>=10'b1001000100) && ({row_reg, col_reg}<10'b1001000110)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}>=10'b1001000110) && ({row_reg, col_reg}<10'b1001001000)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1001001000)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b1001001001)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1001001010)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}>=10'b1001001011) && ({row_reg, col_reg}<10'b1001001111)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1001001111)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1001010000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1001010001)) color_data = 12'b010001000000;
		if(({row_reg, col_reg}==10'b1001010010)) color_data = 12'b010101010000;
		if(({row_reg, col_reg}==10'b1001010011)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1001010100) && ({row_reg, col_reg}<10'b1001011000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1001011000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1001011001) && ({row_reg, col_reg}<10'b1001011011)) color_data = 12'b010101110000;

		if(({row_reg, col_reg}>=10'b1001011011) && ({row_reg, col_reg}<10'b1001100000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1001100000) && ({row_reg, col_reg}<10'b1001100010)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b1001100010)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b1001100011)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1001100100)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}>=10'b1001100101) && ({row_reg, col_reg}<10'b1001101000)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}>=10'b1001101000) && ({row_reg, col_reg}<10'b1001101010)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b1001101010)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}>=10'b1001101011) && ({row_reg, col_reg}<10'b1001110001)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1001110001)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1001110010) && ({row_reg, col_reg}<10'b1001110111)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}>=10'b1001110111) && ({row_reg, col_reg}<10'b1001111001)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1001111001)) color_data = 12'b011110000000;

		if(({row_reg, col_reg}>=10'b1001111010) && ({row_reg, col_reg}<10'b1010000000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1010000000) && ({row_reg, col_reg}<10'b1010000010)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1010000010)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1010000011)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b1010000100)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b1010000101)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1010000110)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}==10'b1010000111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1010001000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b1010001001)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b1010001010)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b1010001011) && ({row_reg, col_reg}<10'b1010001110)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1010001110)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b1010001111)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b1010010000)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b1010010001) && ({row_reg, col_reg}<10'b1010010110)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1010010110)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1010010111)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1010011000) && ({row_reg, col_reg}<10'b1010011100)) color_data = 12'b011110000000;

		if(({row_reg, col_reg}>=10'b1010011100) && ({row_reg, col_reg}<10'b1010100000)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b1010100000) && ({row_reg, col_reg}<10'b1010100010)) color_data = 12'b001101010000;
		if(({row_reg, col_reg}==10'b1010100010)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}==10'b1010100011)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}==10'b1010100100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1010100101)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1010100110)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}==10'b1010100111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1010101000)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b1010101001)) color_data = 12'b100110100001;
		if(({row_reg, col_reg}==10'b1010101010)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}>=10'b1010101011) && ({row_reg, col_reg}<10'b1010101110)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1010101110)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b1010101111) && ({row_reg, col_reg}<10'b1010110010)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b1010110010)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b1010110011)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1010110100)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1010110101)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}>=10'b1010110110) && ({row_reg, col_reg}<10'b1010111000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1010111000) && ({row_reg, col_reg}<10'b1010111010)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1010111010)) color_data = 12'b011110000000;

		if(({row_reg, col_reg}>=10'b1010111011) && ({row_reg, col_reg}<10'b1011000000)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}>=10'b1011000000) && ({row_reg, col_reg}<10'b1011000010)) color_data = 12'b001101010000;
		if(({row_reg, col_reg}==10'b1011000010)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}==10'b1011000011)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b1011000100)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1011000101)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1011000110)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}==10'b1011000111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}>=10'b1011001000) && ({row_reg, col_reg}<10'b1011001010)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1011001010)) color_data = 12'b100110100000;
		if(({row_reg, col_reg}>=10'b1011001011) && ({row_reg, col_reg}<10'b1011001101)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1011001101)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1011001110)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b1011001111) && ({row_reg, col_reg}<10'b1011010010)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b1011010010)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b1011010011)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1011010100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1011010101) && ({row_reg, col_reg}<10'b1011011000)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1011011000)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}==10'b1011011001)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}>=10'b1011011010) && ({row_reg, col_reg}<10'b1011011100)) color_data = 12'b011010000000;

		if(({row_reg, col_reg}>=10'b1011011100) && ({row_reg, col_reg}<10'b1011100000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1011100000)) color_data = 12'b001101010000;
		if(({row_reg, col_reg}==10'b1011100001)) color_data = 12'b001101000000;
		if(({row_reg, col_reg}==10'b1011100010)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}==10'b1011100011)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1011100100)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b1011100101)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1011100110)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}==10'b1011100111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1011101000)) color_data = 12'b101010110001;
		if(({row_reg, col_reg}==10'b1011101001)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1011101010)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b1011101011)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1011101100)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1011101101)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1011101110)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b1011101111) && ({row_reg, col_reg}<10'b1011110001)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b1011110001)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}>=10'b1011110010) && ({row_reg, col_reg}<10'b1011110100)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b1011110100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1011110101)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}>=10'b1011110110) && ({row_reg, col_reg}<10'b1011111010)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1011111010)) color_data = 12'b010001100000;

		if(({row_reg, col_reg}>=10'b1011111011) && ({row_reg, col_reg}<10'b1100000000)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}>=10'b1100000000) && ({row_reg, col_reg}<10'b1100000010)) color_data = 12'b001101010000;
		if(({row_reg, col_reg}==10'b1100000010)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}==10'b1100000011)) color_data = 12'b000000010000;
		if(({row_reg, col_reg}==10'b1100000100)) color_data = 12'b100110110000;
		if(({row_reg, col_reg}==10'b1100000101)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1100000110)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}==10'b1100000111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1100001000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}>=10'b1100001001) && ({row_reg, col_reg}<10'b1100001011)) color_data = 12'b100010100000;
		if(({row_reg, col_reg}==10'b1100001011)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1100001100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1100001101) && ({row_reg, col_reg}<10'b1100010000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1100010000)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b1100010001) && ({row_reg, col_reg}<10'b1100010011)) color_data = 12'b100010010000;
		if(({row_reg, col_reg}==10'b1100010011)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b1100010100)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1100010101)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1100010110) && ({row_reg, col_reg}<10'b1100011000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1100011000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1100011001)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1100011010)) color_data = 12'b010001100000;

		if(({row_reg, col_reg}>=10'b1100011011) && ({row_reg, col_reg}<10'b1100100000)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}==10'b1100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b1100100001) && ({row_reg, col_reg}<10'b1100100011)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}==10'b1100100011)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1100100100)) color_data = 12'b110011010001;
		if(({row_reg, col_reg}>=10'b1100100101) && ({row_reg, col_reg}<10'b1100100111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1100100111)) color_data = 12'b101111000001;
		if(({row_reg, col_reg}==10'b1100101000)) color_data = 12'b100110110001;
		if(({row_reg, col_reg}==10'b1100101001)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}>=10'b1100101010) && ({row_reg, col_reg}<10'b1100101100)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1100101100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1100101101) && ({row_reg, col_reg}<10'b1100101111)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1100101111)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1100110000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1100110001)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b1100110010)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1100110011)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1100110100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1100110101) && ({row_reg, col_reg}<10'b1100111000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1100111000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1100111001)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1100111010)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}==10'b1100111011)) color_data = 12'b001101010000;

		if(({row_reg, col_reg}>=10'b1100111100) && ({row_reg, col_reg}<10'b1101000000)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}>=10'b1101000000) && ({row_reg, col_reg}<10'b1101000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b1101000011) && ({row_reg, col_reg}<10'b1101000111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1101000111)) color_data = 12'b101011000001;
		if(({row_reg, col_reg}==10'b1101001000)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1101001001)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1101001010)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}==10'b1101001011)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1101001100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1101001101)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}>=10'b1101001110) && ({row_reg, col_reg}<10'b1101010000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1101010000)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1101010001)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1101010010)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1101010011)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1101010100)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1101010101) && ({row_reg, col_reg}<10'b1101011001)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1101011001)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1101011010)) color_data = 12'b010001100000;

		if(({row_reg, col_reg}>=10'b1101011011) && ({row_reg, col_reg}<10'b1101100000)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}>=10'b1101100000) && ({row_reg, col_reg}<10'b1101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b1101100011) && ({row_reg, col_reg}<10'b1101101000)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1101101000)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}>=10'b1101101001) && ({row_reg, col_reg}<10'b1101101011)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}>=10'b1101101011) && ({row_reg, col_reg}<10'b1101101111)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1101101111)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1101110000)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1101110001)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1101110010)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1101110011)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1101110100)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1101110101)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}>=10'b1101110110) && ({row_reg, col_reg}<10'b1101111001)) color_data = 12'b011110000000;
		if(({row_reg, col_reg}==10'b1101111001)) color_data = 12'b110011000010;
		if(({row_reg, col_reg}==10'b1101111010)) color_data = 12'b010101110000;

		if(({row_reg, col_reg}>=10'b1101111011) && ({row_reg, col_reg}<10'b1110000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b1110000011) && ({row_reg, col_reg}<10'b1110000110)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1110000110)) color_data = 12'b110011110001;
		if(({row_reg, col_reg}==10'b1110000111)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1110001000)) color_data = 12'b111111110001;
		if(({row_reg, col_reg}>=10'b1110001001) && ({row_reg, col_reg}<10'b1110001011)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}>=10'b1110001011) && ({row_reg, col_reg}<10'b1110001111)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}>=10'b1110001111) && ({row_reg, col_reg}<10'b1110010001)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1110010001)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}==10'b1110010010)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1110010011)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1110010100)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1110010101)) color_data = 12'b100010100001;
		if(({row_reg, col_reg}>=10'b1110010110) && ({row_reg, col_reg}<10'b1110011000)) color_data = 12'b011110000000;

		if(({row_reg, col_reg}>=10'b1110011000) && ({row_reg, col_reg}<10'b1110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=10'b1110100101) && ({row_reg, col_reg}<10'b1110101001)) color_data = 12'b101111010001;
		if(({row_reg, col_reg}==10'b1110101001)) color_data = 12'b011010000000;
		if(({row_reg, col_reg}==10'b1110101010)) color_data = 12'b010001100000;
		if(({row_reg, col_reg}==10'b1110101011)) color_data = 12'b010101010000;
		if(({row_reg, col_reg}>=10'b1110101100) && ({row_reg, col_reg}<10'b1110101110)) color_data = 12'b010101100000;
		if(({row_reg, col_reg}==10'b1110101110)) color_data = 12'b010001010000;
		if(({row_reg, col_reg}==10'b1110101111)) color_data = 12'b010101110000;
		if(({row_reg, col_reg}==10'b1110110000)) color_data = 12'b011001110000;
		if(({row_reg, col_reg}==10'b1110110001)) color_data = 12'b011110010000;
		if(({row_reg, col_reg}>=10'b1110110010) && ({row_reg, col_reg}<10'b1110110100)) color_data = 12'b011110000000;

		if(({row_reg, col_reg}>=10'b1110110100) && ({row_reg, col_reg}<=10'b1110111101)) color_data = 12'b000000000000;
	end
endmodule